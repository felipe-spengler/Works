/*
Usar Clock_25
Contador até 800x525
VGA_HS negativo para H_Sync 660 até 756
Negativo para v 494 até 495
*/
module sign(
	input [11:0]ptx,
	input [11:0]pty,
	input [11:0]p1x,
	input [11:0]p1y,
	input [11:0]p2x,
	input [11:0]p2y,
	output o
	);
	wire signed [11:0] a1;
	wire signed [11:0] a2;
	wire signed [11:0] a3;
	wire signed [11:0] a4;
	wire signed [23:0] m1;
	wire signed [23:0] m2;

	assign a1 = ptx - p2x;
	assign a2 = p1y - p2y;
	assign a3 = p1x - p2x;
	assign a4 = pty - p2y;
	assign m1 = a1 * a2;
	assign m2 = a3 * a4;
	assign o = m1 < m2;

endmodule

module ROM(
	input [4:0]end_triangulo,
	output [11:0]p1x,
	output [11:0]p1y,
	output [11:0]p2x,
	output [11:0]p2y,
	output [11:0]p3x,
	output [11:0]p3y
);

	reg [11:0]p1x_r;
	reg [11:0]p1y_r;
	reg [11:0]p2x_r;
	reg [11:0]p2y_r;
	reg [11:0]p3x_r;
	reg [11:0]p3y_r;

	assign p1x = p1x_r;
	assign p1y = p1y_r;
	assign p2x = p2x_r;
	assign p2y = p2y_r;
	assign p3x = p3x_r;
	assign p3y = p3y_r;

	always @(end_triangulo) begin
		case(end_triangulo)
			0:begin
				p1x_r <= 23;
				p1y_r <= 79;
				p2x_r <= 15;
				p2y_r <= 68;
				p3x_r <= 36;
				p3y_r <= 94;
			end
			1:begin
				p1x_r <= 23;
				p1y_r <= 34;
				p2x_r <= 55;
				p2y_r <= 31;
				p3x_r <= 96;
				p3y_r <= 45;
			end
			2:begin
				p1x_r <= 77;
				p1y_r <= 32;
				p2x_r <= 15;
				p2y_r <= 88;
				p3x_r <= 36;
				p3y_r <= 46;
			end
		endcase
	end
	
endmodule
module video_1(
	input clk,
	input w,
	input [11:0]end_x,
	input [11:0]end_y,
	input data,
	output saida
);
	
	reg memoria_video_1 [0:479] [0:639];
	reg saida_r;
	assign saida = memoria_video_1 [end_x][end_y];
	always @(posedge clk)begin
		if (w == 1) begin
			if (end_x < 640 & end_y < 480)
				memoria_video_1 [end_x][end_y] = data;	
		end	
	end
endmodule
module NewTrab8(
	input CLOCK_50,
	output VGA_HS ,
	output VGA_VS,
	output VGA_R,
	output VGA_G,
	output VGA_B
);
	reg write = 1;

	reg [11:0]p1x;
	reg [11:0]p1y;
	reg [11:0]p2x;
	reg [11:0]p2y;
	reg [11:0]p3x;
	reg [11:0]p3y;
	
	reg [11:0]ptx;
	reg [11:0]pty;

	reg [11:0]i;
	reg [11:0]j;
	
	wire [11:0]ptx_w;
	wire [11:0]pty_w;
	wire [11:0]p1x_w;
	wire [11:0]p1y_w;
	wire [11:0]p2x_w;
	wire [11:0]p2y_w;
	wire [11:0]p3x_w;
	wire [11:0]p3y_w;	

	reg [3:0]count = 0;
	reg [4:0]end_triangulo = 0;
	wire P1, P2, P3;
	reg saida;
	wire data;

	reg pode_ler = 0;
	
	reg [3:0]Red;
	reg [3:0]Green;
	reg [3:0]Blue;
	reg [11:0]V_Sync;
	reg [11:0]H_Sync;

	reg CLK_25 = 0;

	assign VGA_R = Red;
	assign VGA_B = Blue;
	assign VGA_G = Green;
	
	assign VGA_HS = H_Sync;
	assign VGA_VS = V_Sync;
	
	sign Pt1(ptx, pty, p1x, p1y, p2x, p2y, P1);
	sign Pt2(ptx, pty, p2x, p2y, p3x, p3y, P2);
	sign Pt3(ptx, pty, p3x, p3y, p1x, p1y, P3);
	ROM R(end_triangulo, p1x_w, p1y_w, p2x_w, p2y_w, p3x_w, p3y_w);
	video_1 V(CLK_25, write, i, j, saida, data); 

	always @(posedge CLOCK_50) CLK_25 <= ~CLK_25;
	always @(posedge CLK_25) begin
		case(count)
			0:begin
				end_triangulo <= 0;
				count <= 1;
			end
			1: begin
				$display (" Triangulo %d", end_triangulo);
				p1x <= p1x_w;
				p1y <= p1y_w;
				p2x <= p2x_w;
				p2y <= p2y_w;
				p3x <= p3x_w;
				p3y <= p3y_w;	

				i <= 0;
				j <= 0;
				count <= 2;
				if (end_triangulo > 2) write <= 0;
				else write <= 1;
			end

			
			2: begin
				if (i < 640)begin
					count <= 3;
					j <= 0;
					
				end
		    		else count <= 4;
			end
			3: begin
				if (j < 480)begin
					// sempe alterar aqui (dentro for)
					ptx <= i;
					pty <= j;
					
					if (i  > 660 & i < 756) H_Sync <= 0;
					else H_Sync <= 1;
               if (j  > 494 & j < 495) V_Sync <= 0;
					else V_Sync <= 1;
					
					saida <= P1 == P2 & P2 == P3;

					if (pode_ler == 1)begin
						
						if (data == 1)begin
							Red <= 4'b1;
							Green <= 4'b1;
							Blue <= 4'b1;
						end
						else begin
							Red <= 4'b0;
							Green <= 4'b0;
							Blue <= 4'b0;
						end
					end
					//altera até aqui (dentro for)
					j <= j + 1;
					count <= 3;	
				end
				else begin
					i <= i + 1;
					count = 2;
				end
			end
			4: begin
				count <= 5;
				write <= 0;
			end


			5: begin
				if (pode_ler == 0) pode_ler <= 1;
				end_triangulo <= end_triangulo + 1;
				count <= 6;
			end
			6:begin
				if (end_triangulo > 3) $finish;
				else count <= 1;
			end
			
		endcase
	end	

endmodule

